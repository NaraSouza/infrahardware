module mux_pccond(
	//TODO: Verificar se output est� correto
	input wire [1:0] selector,
	input wire equal,//00
	input wire greater,//01
	output wire out);
	
	
always
	case(selector)
		2'b00: out = equal;
		2'b01: out = !equal;
		2'b10: out = !greater;
		2'b11: out = greater;
endcase
	
endmodule: mux_pccond