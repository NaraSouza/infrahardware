module CPU(input clock,
	input reset,
	output logic [31:0] pcout,
	output logic [31:0] epcout,
	output logic [31:0] mdrout,
	output logic [5:0] op,
	output logic [4:0] rs,
    output logic [4:0] rt,
    output logic [15:0] inst15_0,
	output logic [6:0] stateout
);

//fios grandoes:
logic pccontrol;
logic [31:0] wmwritedata;
logic [31:0] alusrcaout;
logic [31:0] alusrcbout;
logic [31:0] regaluout;
logic [31:0] memtoregout;
logic [2:0] aluop;
logic [31:0] regdeslocout;
logic memwrite;
logic regwritesignal;
logic irwrite;
logic [31:0] regaout;
logic [31:0] regbout;
logic [4:0] shamt;
logic [2:0] shiftop;
logic [4:0] regdstout;
logic [1:0] readdstmux;
logic readsmux;
logic [31:0] regain;
logic [4:0] shiftsout;
logic [31:0] reginout;
logic [31:0] aluresult;
logic [31:0] highout;
logic [31:0] lowout;	
logic [31:0] iordout;



logic pcond1;
logic ltflag;
logic equalflag;
logic gtflag;
logic pccond2;
logic [5:0] funct;
logic [31:0] memout;
logic [31:0] pcin;
logic [31:0] wmregout;
logic [25:0] inst25_0; //facilita ter s� ele porque no 
 //n�o precisa concatenar nada
logic [4:0] rd;
logic [4:0] sp; //$29
logic [4:0] reg31; //$31
logic [4:0] readsout; 
logic [31:0] signextendout;
logic [31:0] sl1out;
logic [31:0] sl2out;
logic [31:0] regbin;

logic [31:0] divhighout;
logic [31:0] divlowout;
logic [31:0] multhighout;
logic [31:0] multlowout;
logic [31:0] muxhighout;
logic [31:0] muxlowout;
logic [31:0] multsout;

//sinais de pc:
logic pccondout; //saida do mux pccond
logic pcwritecond; // sinal da unidade de controle
logic pcwrite; // sinal da unidade de controle
logic pcand; //pcwritecond and pccondout
 //fio da unidade de controle que entra em pc (pcand or pcwrite)

assign pcand = pcwritecond && pccondout;
assign pccontrol = pcand || pcwrite;

//sinais de registradores:
logic mdrs;
logic regaw;
logic regbw;
logic regaluwrite;
logic epcwrite;
logic reghighw;
logic regloww;

//sinais dos mux:
logic [2:0] iordmux; //mux 5 //mux 2 //mux 4
logic [2:0] memtoregmux; //mux 7
logic alusrcamux; //mux 2
logic [1:0] alusrcbmux; //mux 4
logic [2:0] pcsourcemux; //mux 6
logic reginmux; //mux 2
logic shiftsmux; //mux 2
logic divmultmux; //mux 2
logic multsmux; //mux 2
logic [1:0] pccondmux;

// sinais dos componentes:
logic [1:0] wms; //write mode signal

logic startdiv;
logic divstop;
logic divzero;
logic startmult;
logic stopmult;
logic multo;

// saidas da ula:
logic zeroflag;
logic negflag;
logic overflowflag;



endmodule: CPU